`ifndef _s32
`define _s32
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date:    16:36:55 11/15/2017
// Design Name:
// Module Name:    Shift32
// Project Name:
// Target Devices:
// Tool versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
module Shift32(in, out);

	input [31:0] in;
	output [31:0] out;
	assign out = in << 2;

endmodule
`endif
